module and2
(
	input a, 
	input b, 
	output andOut
);

assign andOut = a & b;

endmodule