4x4 Multiplier 

.include TSMC_180nm.txt
.param w=360n
.param l=180n
.param vdd_val=0.8
VDD Vdd GND vdd_val 

*subckts*

.SUBCKT AND input1_and input2_and output Vdd
Mp1 node1_AND    input1_and       Vdd Vdd CMOSP W={w} L=l
Mp2 node1_AND    input2_and       Vdd Vdd CMOSP W={w} L=l
Mp3    output     node1_AND       Vdd Vdd CMOSP   W=w L=l
Mn1 node1_AND    input1_and node2_AND GND CMOSN W={w} L=l
Mn2 node2_AND    input2_and       GND GND CMOSN W={w} L=l
Mn3    output     node1_AND       GND GND CMOSN W={2*w} L=l
.ENDS AND 

.SUBCKT FULL_ADDER input1 input2 input3 sum carry Vdd 
 Mp1  node1 input1    Vdd Vdd CMOSP    W={2*w} L=l
 Mp2  node2 input2  node1 Vdd CMOSP    W={2*w} L=l
 Mp3  node4 input1    Vdd Vdd CMOSP    W={2*w} L=l
 Mp4  node4 input2    Vdd Vdd CMOSP    W={2*w} L=l
 Mp5  node2 input3  node4 Vdd CMOSP    W={2*w} L=l
 Mp6  node6 input3    Vdd Vdd CMOSP    W={2*w} L=l
 Mp7  node6 input2    Vdd Vdd CMOSP    W={2*w} L=l
 Mp8  node6 input1    Vdd Vdd CMOSP    W={2*w} L=l
 Mp9  node8  node2  node6 Vdd CMOSP    W={2*w} L=l
Mp10  node9 input1    Vdd Vdd CMOSP W={1.33*w} L=l
Mp11 node10 input2  node9 Vdd CMOSP W={1.33*w} L=l
Mp12  node8 input3 node10 Vdd CMOSP W={1.33*w} L=l
Mp13    sum  node8    Vdd Vdd CMOSP    W={4*w} L=l
Mp14  carry  node2    Vdd Vdd CMOSP    W={4*w} L=l
 Mn1  node2 input2  node3 GND CMOSN        W=w L=l
 Mn2  node3 input1    GND GND CMOSN        W=w L=l
 Mn3  node2 input3  node5 GND CMOSN        W=w L=l
 Mn4  node5 input1    GND GND CMOSN        W=w L=l
 Mn5  node5 input2    GND GND CMOSN        W=w L=l
 Mn6  node8  node2  node7 GND CMOSN        W=w L=l
 Mn7  node7 input3    GND GND CMOSN        W=w L=l
 Mn8  node7 input2    GND GND CMOSN        W=w L=l
 Mn9  node7 input1    GND GND CMOSN        W=w L=l
Mn10  node8 input3 node11 GND CMOSN W={0.66*w} L=l
Mn11 node11 input2 node12 GND CMOSN W={0.66*w} L=l
Mn12 node12 input1    GND GND CMOSN W={0.66*w} L=l
Mn13    sum  node8    GND GND CMOSN    W={2*w} L=l
MN14  carry  node2    GND GND CMOSN    W={2*w} L=l
.ENDS FULL_ADDER

.SUBCKT HALF_ADDER input1_half input2_half sum_half carry_half Vdd
Mp1    node1_half       node9_half        Vdd Vdd CMOSP W={2*w} L=l
Mp2  	 sum_half      input2_half node1_half Vdd CMOSP W={2*w} L=l
Mp3    node2_half      input1_half        Vdd Vdd CMOSP W={2*w} L=l
Mp4 	 sum_half       node8_half node2_half Vdd CMOSP W={2*w} L=l
Mp5    node6_half  	node9_half        Vdd Vdd CMOSP W={2*w} L=l
Mp6    carry_half  	node8_half node6_half Vdd CMOSP W={2*w} L=l
Mp7    node8_half      input2_half        Vdd Vdd CMOSP W={4*w} L=l
Mp8    node9_half      input1_half        Vdd Vdd CMOSP W={4*w} L=l
Mn1 	 sum_half      input1_half node4_half GND CMOSN     W=w L=l
Mn2    node4_half      input2_half        GND GND CMOSN     W=w L=l
Mn3 	 sum_half  	node9_half node5_half GND CMOSN     W=w L=l
Mn4    node5_half  	node8_half        GND GND CMOSN     W=w L=l
Mn5    carry_half  	node9_half        GND GND CMOSN W={4*w} L=l
Mn6    carry_half  	node8_half        GND GND CMOSN W={4*w} L=l
Mn7    node8_half      input2_half        GND GND CMOSN W={4*w} L=l
Mn8    node9_half      input1_half        GND GND CMOSN W={4*w} L=l
.ENDS HALF_ADDER

 X1  input1    input5   P0  Vdd  		AND
 X2  input2    input5   K2  Vdd  		AND
 X3  input3    input5   K3  Vdd  		AND
 X4  input4    input5   K4  Vdd  		AND
 X5  input1    input6   K5  Vdd  		AND
 X6  input2    input6   K6  Vdd  		AND
 X7  input3    input6   K7  Vdd  		AND
 X8  input4    input6   K8  Vdd  		AND
 X9      K5        K2   P1 CHA1  Vdd 	 HALF_ADDER
X10      K6        K3 CHA1 SFA1 CFA1 Vdd FULL_ADDER
X11      K7        K4 CFA1 SFA2 CFA2 Vdd FULL_ADDER
X12      K8      CFA2 SHA2 CHA2  Vdd 	 HALF_ADDER
X13  input1    input7   K9  Vdd  		AND
X14  input2    input7  K10  Vdd  		AND
X15  input3    input7  K11  Vdd  		AND
X16  input4    input7  K12  Vdd                 AND
X17      K9      SFA1   P2 CHA3  Vdd 	 HALF_ADDER
X18    CHA3       K10 SFA2 SFA3 CFA3 Vdd FULL_ADDER
X19     K11      CFA3 SHA2 SFA4 CFA4 Vdd FULL_ADDER
X20     K12      CFA4 CHA2 SFA5 CFA5 Vdd FULL_ADDER
X21  input1    input8  K13  Vdd 		AND
X22  input2    input8  K14  Vdd 		AND
X23  input3    input8  K15  Vdd 		AND
X24  input4    input8  K16  Vdd 		AND
X25     K13      SFA3   P3 CHA4  Vdd 	 HALF_ADDER
X26     K14      CHA4 SFA4   P4 CFA6 Vdd FULL_ADDER
X27     K15      CFA6 SFA5   P5 CFA7 Vdd FULL_ADDER
X28     K16      CFA7 CFA5   P6   P7 Vdd FULL_ADDER 

Cp0 P0 GND 1.0f
Cp1 P1 GND 1.0f
Cp2 P2 GND 1.0f
Cp3 P3 GND 1.0f
Cp4 P4 GND 1.0f
Cp5 P5 GND 1.0f
Cp6 P6 GND 1.0f
Cp7 P7 GND 1.0f

V7 input8 0 DC=0 PULSE(0 vdd_val 3200u 100n 100n 3200u  6400u)
V6 input7 0 DC=0 PULSE(0 vdd_val 1600u 100n 100n 1600u  3200u)
V5 input6 0 DC=0 PULSE(0 vdd_val  800u 100n 100n  800u  1600u)
V4 input5 0 DC=0 PULSE(0 vdd_val  400u 100n 100n  400u   800u)
V3 input4 0 DC=0 PULSE(0 vdd_val  200u 100n 100n  200u   400u)
V2 input3 0 DC=0 PULSE(0 vdd_val  100u 100n 100n  100u   200u)
V1 input2 0 DC=0 PULSE(0 vdd_val   50u 100n 100n   50u   100u)
V0 input1 0 DC=0 PULSE(0 vdd_val   25u 100n 100n   25u    50u) 

.control
tran 25us 12456us 10us 

let delay_LH_P6 = 0
let delay_HL_P6 = 0

meas tran delay_LH_P6 trig v(input2) val = 0.5 rise = 31 targ v(P6) val = 0.5 rise = 10
meas tran delay_HL_P6 trig v(input2) val = 0.5 fall = 24 targ v(P6) val = 0.5  fall = 5

let avg_delay_P6 = (delay_LH_P6 + delay_HL_P6)/2

echo                           " ---------------------------------------"  > "multiplier_delays.txt"
echo "|-> low to high delay worst case = "               "$&delay_LH_P6|" >> "multiplier_delays.txt"
echo "|-> high to low delay worst case = "          "     $&delay_HL_P6|" >> "multiplier_delays.txt"
echo "|->  worst case delay (P6) = " 	           "     $&avg_delay_P6|" >> "multiplier_delays.txt"
echo                           " ---------------------------------------" >> "multiplier_delays.txt"

.endc
.end

