FULL ADDER

.include TSMC_180nm.txt
.param w=360n
.param l=180n
.param vdd_val=1
*********
*Netlist*
*********

VDD Vdd GND vdd_val

*mos D G S B model W L
 Mp1  node1 input1    Vdd Vdd CMOSP    W={2*w} L=l
 Mp2  node2 input2  node1 Vdd CMOSP    W={2*w} L=l
 Mp3  node4 input1    Vdd Vdd CMOSP    W={2*w} L=l
 Mp4  node4 input2    Vdd Vdd CMOSP    W={2*w} L=l
 Mp5  node2 input3  node4 Vdd CMOSP    W={2*w} L=l
 Mp6  node6 input3    Vdd Vdd CMOSP    W={2*w} L=l
 Mp7  node6 input2    Vdd Vdd CMOSP    W={2*w} L=l
 Mp8  node6 input1    Vdd Vdd CMOSP    W={2*w} L=l
 Mp9  node8  node2  node6 Vdd CMOSP    W={2*w} L=l
Mp10  node9 input1    Vdd Vdd CMOSP W={1.33*w} L=l
Mp11 node10 input2  node9 Vdd CMOSP W={1.33*w} L=l
Mp12  node8 input3 node10 Vdd CMOSP W={1.33*w} L=l
Mp13    sum  node8    Vdd Vdd CMOSP    W={4*w} L=l
Mp14  carry  node2    Vdd Vdd CMOSP    W={4*w} L=l
 Mn1  node2 input2  node3 GND CMOSN        W=w L=l
 Mn2  node3 input1    GND GND CMOSN        W=w L=l
 Mn3  node2 input3  node5 GND CMOSN        W=w L=l
 Mn4  node5 input1    GND GND CMOSN        W=w L=l
 Mn5  node5 input2    GND GND CMOSN        W=w L=l
 Mn6  node8  node2  node7 GND CMOSN        W=w L=l
 Mn7  node7 input3    GND GND CMOSN        W=w L=l
 Mn8  node7 input2    GND GND CMOSN        W=w L=l
 Mn9  node7 input1    GND GND CMOSN        W=w L=l
Mn10  node8 input3 node11 GND CMOSN W={0.66*w} L=l
Mn11 node11 input2 node12 GND CMOSN W={0.66*w} L=l
Mn12 node12 input1    GND GND CMOSN W={0.66*w} L=l
Mn13    sum  node8    GND GND CMOSN    W={2*w} L=l
MN14  carry  node2    GND GND CMOSN    W={2*w} L=l

CoutS   sum GND 1.5f
CoutC carry GND 1.5f

V2 input3 0 DC=0 PULSE(0 vdd_val 200u 100n 100n 200u 400u)
V1 input2 0 DC=0 PULSE(0 vdd_val 100u 100n 100n 100u 200u)
V0 input1 0 DC=0 PULSE(0 vdd_val  50u 100n 100n  50u 100u)

*control*

.control

tran 25us 1625us 

plot v(input1) 
plot v(input2)
plot v(input3)
plot    v(sum)
plot  v(carry)

let delay_sum_LH = 0
let delay_sum_HL = 0
let delay_carry_LH = 0
let delay_carry_HL = 0
meas tran   delay_sum_LH trig v(input1) val = 0.5 rise = 1 targ   v(sum) val = 0.5 rise = 1
meas tran   delay_sum_HL trig v(input1) val = 0.5 rise = 2 targ   v(sum) val = 0.5 fall = 2
meas tran delay_carry_LH trig v(input1) val = 0.5 rise = 2 targ v(carry) val = 0.5 rise = 2
meas tran delay_carry_HL trig v(input1) val = 0.5 fall = 4 targ v(carry) val = 0.5 fall = 3

let propDelSum = (abs(delay_sum_LH) + abs(delay_sum_HL))/2
let propDelcarry = (abs(delay_carry_LH) + abs(delay_carry_HL))/2
echo				  " -----------------------------------------------------------" > "output_full_adder.txt"
echo 	"|->            high to low delay_sum = " 	"		     $&delay_sum_HL|"   >> "output_full_adder.txt"
echo "|-> 	       low to high delay_sum = " 	  "	       $&delay_sum_LH|"         >> "output_full_adder.txt"
echo 		"|-> worst case propogation delay_sum = " "		$&propDelSum|"          >> "output_full_adder.txt"
echo " -----------------------------------------------------------" >> "output_full_adder.txt"
echo   "|->            high to low delay_carry = " 	"		     $&delay_carry_HL|" >> "output_full_adder.txt"
echo "|-> 	       low to high delay_carry = " 	"	       $&delay_carry_LH|"       >> "output_full_adder.txt"
echo   "|-> worst case propogation delay_carry = " 	"		$&propDelcarry|"        >> "output_full_adder.txt"
echo 				 " -----------------------------------------------------------" >> "output_full_adder.txt"


.endc
.end
