AND gate 

.include TSMC_180nm.txt
.param w=360n 
.param l=180n
.param vdd_val=1

*********
*Netlist*
*********

VDD vdd GND vdd_val

*mos D G S B model W L

Mp1 node1 nodeA   vdd vdd CMOSP   W={w} L=l
Mp2 node1 nodeB   vdd vdd CMOSP   W={w} L=l
Mp3   out node1   vdd vdd CMOSP   W={w} L=l
Mn1 node1 nodeA node2 GND CMOSN   W={w} L=l
Mn2 node2 nodeB   GND GND CMOSN   W={w} L=l
Mn3   out node1   GND GND CMOSN W={2*w} L=l

Cout out GND 1.5f

Va nodeA GND pulse(0 vdd_val 0 0.1n 0.1n 10n 20n)
Vb nodeB GND pulse(0 vdd_val 0 0.1n 0.1n 20n 40n)

.control
tran 0.1n 100n

plot   v(out) 
plot v(nodeA)
plot v(nodeB)

let delay_and_lh = 0
let delay_and_hl = 0

meas tran delay_and_lh trig v(nodeA) val = 0.5 rise = 1 targ v(out) val = 0.5 rise = 1
meas tran delay_and_hl trig v(nodeA) val = 0.5 fall = 1 targ v(out) val = 0.5 fall = 1
let prop_del_and = (delay_and_lh + delay_and_hl)/2

echo                                              " ---------------------------------"  > "and_delays.txt"
echo 					  "|-> low to high delay = " "$&delay_and_lh|" >> "and_delays.txt"
echo 					  "|-> high to low delay = " "$&delay_and_hl|" >> "and_delays.txt"
echo 			          "|-> average propogation delay = " "$&prop_del_and|" >> "and_delays.txt"
echo                            	          " ---------------------------------" >> "and_delays.txt"

.endc
.end
