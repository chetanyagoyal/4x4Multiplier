HALF ADDER 

.include TSMC_180nm.txt
.param w=360n
.param l=180n
.param vdd_val=1

*********
*Netlist*
*********

VDD vdd GND vdd_val

*mos D G S B model W L

Mp1    node1_half       node9_half        Vdd Vdd CMOSP W={2*w} L=l
Mp2  	 sum_half      input2_half node1_half Vdd CMOSP W={2*w} L=l
Mp3    node2_half      input1_half        Vdd Vdd CMOSP W={2*w} L=l
Mp4 	 sum_half       node8_half node2_half Vdd CMOSP W={2*w} L=l
Mp5    node6_half  	node9_half        Vdd Vdd CMOSP W={2*w} L=l
Mp6    carry_half  	node8_half node6_half Vdd CMOSP W={2*w} L=l
Mp7    node8_half      input2_half        Vdd Vdd CMOSP W={4*w} L=l
Mp8    node9_half      input1_half        Vdd Vdd CMOSP W={4*w} L=l
Mn1 	 sum_half      input1_half node4_half GND CMOSN     W=w L=l
Mn2    node4_half      input2_half        GND GND CMOSN     W=w L=l
Mn3 	 sum_half  	node9_half node5_half GND CMOSN     W=w L=l
Mn4    node5_half  	node8_half        GND GND CMOSN     W=w L=l
Mn5    carry_half  	node9_half        GND GND CMOSN W={4*w} L=l
Mn6    carry_half  	node8_half        GND GND CMOSN W={4*w} L=l
Mn7    node8_half      input2_half        GND GND CMOSN W={4*w} L=l
Mn8    node9_half      input1_half        GND GND CMOSN W={4*w} L=l

CoutS   sum_half GND 1.5f
CoutC carry_half GND 1.5f

V1 input2_half 0 DC=0 PULSE(0 vdd_val  100u 100n 100n  100u   200u)
V0 input1_half 0 DC=0 PULSE(0 vdd_val   50u 100n 100n   50u   100u)

*control*
.control 

tran 25us 1625us

plot v(sum_half) 
plot v(input2_half) 
plot v(input1_half)
plot v(carry_half)

let delay_in1_LH = 0
let delay_carry_LH = 0
let delay_in1_HL = 0
let delay_carry_HL = 0
meas tran delay_in1_LH trig v(input1_half) val = 0.5 rise = 3 targ v(sum_half) val = 0.5 rise = 3
meas tran delay_in1_HL trig v(input1_half) val = 0.5 rise = 2 targ v(sum_half) val = 0.5 fall = 2
meas tran delay_carry_LH trig v(input1_half) val = 0.5 rise = 2 targ v(carry_half) val = 0.5 rise = 2
meas tran delay_carry_HL trig v(input1_half) val = 0.5 fall = 6 targ v(carry_half) val = 0.5 fall = 6
let   propDelIn1 =          (abs(delay_in1_LH) + abs(delay_in1_HL))/2
let propDelcarry = 	(abs(delay_carry_LH) + abs(delay_carry_HL))/2

echo " ---------------------------------------------"                 > "output_half_adder.txt"
echo "|->            low to high delay_sum = " "$&delay_in1_LH|"     >> "output_half_adder.txt"
echo "|->            high to low delay_sum = " "$&delay_in1_HL|"     >> "output_half_adder.txt"
echo "|-> worst case propogation delay_sum = " " $&propDelIn1|"      >> "output_half_adder.txt"
echo " ---------------------------------------------"		     >> "output_half_adder.txt"
echo " ---------------------------------------------" 		     >> "output_half_adder.txt"
echo "|->            low to high delay_carry = " "$&delay_carry_LH|" >> "output_half_adder.txt"
echo "|->            high to low delay_carry = " "$&delay_carry_HL|" >> "output_half_adder.txt"
echo "|-> worst case propogation delay_carry = " " $&propDelcarry|"  >> "output_half_adder.txt"
echo " ---------------------------------------------"                >> "output_half_adder.txt"
.endc
.end
