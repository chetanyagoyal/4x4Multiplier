magic
tech scmos
timestamp 1669480491
<< nwell >>
rect -6 -6 47 23
rect 54 -3 100 24
<< ntransistor >>
rect 8 -27 12 -19
rect 29 -27 33 -19
rect 75 -23 79 -19
<< ptransistor >>
rect 8 0 12 8
rect 29 0 33 8
rect 75 3 79 11
<< ndiffusion >>
rect 7 -27 8 -19
rect 12 -27 29 -19
rect 33 -27 34 -19
rect 65 -23 75 -19
rect 79 -23 88 -19
<< pdiffusion >>
rect 7 0 8 8
rect 12 0 17 8
rect 24 0 29 8
rect 33 0 34 8
rect 65 3 75 11
rect 79 3 88 11
<< ndcontact >>
rect 0 -27 7 -19
rect 34 -27 41 -19
rect 60 -23 65 -19
rect 88 -23 93 -19
<< pdcontact >>
rect 0 0 7 8
rect 17 0 24 8
rect 34 0 41 8
rect 60 3 65 11
rect 88 3 93 11
<< psubstratepcontact >>
rect 0 -38 7 -32
rect 60 -38 65 -32
<< nsubstratencontact >>
rect 0 13 7 18
rect 34 13 41 18
rect 60 15 65 19
<< polysilicon >>
rect 8 8 12 17
rect 29 8 33 17
rect 75 11 79 15
rect 8 -19 12 0
rect 29 -19 33 0
rect 75 -19 79 3
rect 75 -26 79 -23
rect 8 -30 12 -27
rect 29 -30 33 -27
<< polycontact >>
rect 70 -15 75 -10
<< metal1 >>
rect 0 19 65 25
rect 0 18 7 19
rect 0 8 7 13
rect 34 18 41 19
rect 34 8 41 13
rect 60 11 65 15
rect 17 -10 24 0
rect 17 -15 70 -10
rect 34 -19 41 -15
rect 88 -19 93 3
rect 0 -32 7 -27
rect 60 -32 65 -23
rect 7 -38 60 -32
<< end >>
