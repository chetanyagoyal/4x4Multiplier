magic
tech scmos
timestamp 1669569837
<< nwell >>
rect 0 0 59 47
rect 70 0 129 48
rect 0 -116 41 -86
rect 67 -112 108 -91
rect 5 -173 63 -145
rect 71 -176 112 -151
<< ntransistor >>
rect 15 -40 19 -32
rect 40 -40 44 -32
rect 85 -40 89 -32
rect 110 -40 114 -32
rect 18 -78 22 -74
rect 85 -84 89 -80
rect 18 -198 22 -182
rect 46 -198 50 -182
rect 89 -188 93 -184
<< ptransistor >>
rect 15 7 19 23
rect 40 7 44 23
rect 85 7 89 23
rect 110 7 114 23
rect 18 -100 22 -92
rect 85 -105 89 -97
rect 18 -167 22 -159
rect 46 -167 50 -159
rect 89 -170 93 -162
<< ndiffusion >>
rect 14 -40 15 -32
rect 19 -40 40 -32
rect 44 -40 45 -32
rect 84 -40 85 -32
rect 89 -40 110 -32
rect 114 -40 115 -32
rect 11 -78 18 -74
rect 22 -78 30 -74
rect 78 -84 85 -80
rect 89 -84 97 -80
rect 17 -198 18 -182
rect 22 -198 46 -182
rect 50 -198 51 -182
rect 82 -188 89 -184
rect 93 -188 101 -184
<< pdiffusion >>
rect 14 7 15 23
rect 19 7 40 23
rect 44 7 45 23
rect 84 7 85 23
rect 89 7 110 23
rect 114 7 115 23
rect 11 -100 18 -92
rect 22 -100 30 -92
rect 78 -105 85 -97
rect 89 -105 97 -97
rect 17 -167 18 -159
rect 22 -167 31 -159
rect 37 -167 46 -159
rect 50 -167 51 -159
rect 82 -170 89 -162
rect 93 -170 101 -162
<< ndcontact >>
rect 6 -40 14 -32
rect 45 -40 53 -32
rect 76 -40 84 -32
rect 115 -40 123 -32
rect 6 -78 11 -74
rect 30 -78 35 -74
rect 73 -84 78 -80
rect 97 -84 102 -80
rect 11 -198 17 -182
rect 51 -198 57 -182
rect 77 -188 82 -184
rect 101 -188 106 -184
<< pdcontact >>
rect 6 7 14 23
rect 45 7 53 23
rect 76 7 84 23
rect 115 7 123 23
rect 6 -100 11 -92
rect 30 -100 35 -92
rect 73 -105 78 -97
rect 97 -105 102 -97
rect 11 -167 17 -159
rect 31 -167 37 -159
rect 51 -167 57 -159
rect 77 -170 82 -162
rect 101 -170 106 -162
<< psubstratepcontact >>
rect 6 -50 14 -44
rect 6 -70 11 -66
rect 76 -50 84 -45
rect 73 -76 78 -72
rect 77 -197 82 -192
rect 11 -207 17 -202
<< nsubstratencontact >>
rect 6 36 14 42
rect 76 36 84 42
rect 6 -113 11 -108
rect 11 -152 17 -148
rect 73 -123 78 -118
rect 51 -153 57 -148
rect 77 -158 82 -154
<< polysilicon >>
rect 15 44 137 48
rect 15 23 19 44
rect 40 23 44 34
rect 85 23 89 35
rect 110 23 114 34
rect 15 -3 19 7
rect 40 -18 44 7
rect 85 -1 89 7
rect 15 -22 44 -18
rect 69 -5 89 -1
rect 15 -32 19 -22
rect 40 -32 44 -26
rect 15 -56 19 -40
rect 40 -44 44 -40
rect 69 -44 73 -5
rect 110 -9 114 7
rect 85 -13 114 -9
rect 85 -32 89 -13
rect 110 -32 114 -29
rect 40 -48 73 -44
rect 15 -60 22 -56
rect 18 -74 22 -60
rect 69 -67 73 -48
rect 85 -57 89 -40
rect 110 -43 114 -40
rect 133 -43 137 44
rect 114 -47 137 -43
rect 69 -71 89 -67
rect 18 -92 22 -78
rect 85 -80 89 -71
rect 85 -97 89 -84
rect 18 -159 22 -100
rect 85 -113 89 -105
rect 46 -117 89 -113
rect 46 -159 50 -117
rect 89 -162 93 -151
rect 18 -182 22 -167
rect 46 -182 50 -167
rect 89 -184 93 -170
rect 89 -192 93 -188
rect 18 -201 22 -198
rect 46 -201 50 -198
<< polycontact >>
rect 110 -47 114 -43
rect 85 -62 89 -57
rect 84 -181 89 -177
<< metal1 >>
rect 14 36 76 42
rect 84 36 145 42
rect 6 23 14 36
rect 76 23 84 36
rect 45 -10 53 7
rect 115 -10 123 7
rect 45 -17 123 -10
rect 45 -32 53 -17
rect 57 -28 102 -23
rect 6 -44 14 -40
rect 57 -49 62 -28
rect 76 -45 84 -40
rect 14 -50 76 -49
rect 6 -54 84 -50
rect 6 -62 11 -54
rect -11 -66 11 -62
rect 85 -64 89 -62
rect -11 -67 6 -66
rect -11 -111 -5 -67
rect 6 -74 11 -70
rect 42 -68 89 -64
rect 30 -80 35 -78
rect 42 -80 47 -68
rect 98 -71 102 -28
rect 115 -32 123 -17
rect 30 -84 47 -80
rect 73 -72 102 -71
rect 78 -75 102 -72
rect 73 -80 78 -76
rect 30 -92 35 -84
rect 97 -85 102 -84
rect 110 -85 114 -47
rect 139 -50 145 36
rect 97 -89 114 -85
rect 118 -55 145 -50
rect 97 -97 102 -89
rect 6 -108 11 -100
rect -11 -116 2 -111
rect -4 -207 2 -116
rect 6 -118 11 -113
rect 73 -118 78 -105
rect 118 -118 124 -55
rect 6 -123 73 -118
rect 78 -123 124 -118
rect 33 -131 38 -123
rect 11 -136 82 -131
rect 11 -148 17 -136
rect 11 -159 17 -152
rect 51 -148 57 -136
rect 51 -159 57 -153
rect 77 -154 82 -136
rect 77 -162 82 -158
rect 31 -177 37 -167
rect 31 -181 84 -177
rect 101 -178 106 -170
rect 51 -182 57 -181
rect 101 -182 118 -178
rect 101 -184 106 -182
rect 77 -192 82 -188
rect 11 -202 17 -198
rect 77 -207 82 -197
rect -4 -212 82 -207
<< end >>
