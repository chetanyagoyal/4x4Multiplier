magic
tech scmos
timestamp 1669380902
<< polysilicon >>
rect 0 105 240 109
rect 0 92 4 105
rect 79 92 83 105
rect 162 92 166 105
rect 236 92 240 105
rect 8 76 314 80
rect -7 55 10 59
rect 75 55 89 59
rect 159 55 172 59
rect 231 55 245 59
rect 287 55 364 59
rect -7 17 -3 55
rect -25 13 -3 17
rect -606 -242 -601 -94
rect -25 -100 -21 13
rect -7 -31 -3 13
rect 57 -18 61 23
rect 71 -31 75 55
rect 138 -2 142 23
rect 138 -6 147 -2
rect 143 -18 147 -6
rect 155 -31 159 55
rect 221 -5 225 23
rect 231 3 235 55
rect 231 -1 242 3
rect 221 -9 231 -5
rect 227 -18 231 -9
rect 238 -31 242 -1
rect 295 -5 299 23
rect 295 -9 311 -5
rect 307 -18 311 -9
rect -7 -35 7 -31
rect 71 -35 92 -31
rect 155 -35 176 -31
rect 238 -35 257 -31
rect 52 -56 93 -52
rect 139 -56 176 -52
rect 223 -56 260 -52
rect 303 -56 318 -52
rect -441 -104 -21 -100
rect -522 -161 -518 -125
rect -509 -157 -505 -137
rect -509 -160 -490 -157
rect -445 -523 -441 -104
rect -434 -116 -430 -114
rect -434 -120 -137 -116
rect -434 -366 -430 -120
rect -141 -158 -137 -120
rect -221 -333 -149 -329
rect -426 -344 -418 -339
rect -434 -370 -414 -366
rect -445 -527 -258 -523
rect -262 -612 -258 -527
rect -262 -616 -204 -612
rect -208 -664 -204 -616
rect -132 -664 -128 -113
rect 57 -115 61 -88
rect 143 -115 147 -88
rect 227 -115 231 -88
rect 307 -115 311 -88
rect 360 -110 364 55
rect 360 -114 396 -110
rect 57 -119 311 -115
rect 57 -144 61 -119
rect -115 -148 61 -144
rect -115 -154 -111 -148
rect 225 -232 229 -119
rect 299 -160 303 -143
rect 317 -157 321 -142
rect 317 -161 331 -157
rect -108 -356 -47 -352
rect -123 -635 -119 -503
rect -108 -537 -104 -356
rect 392 -431 396 -114
rect 212 -435 396 -431
rect -108 -541 41 -537
rect -691 -668 -104 -664
rect -783 -692 -440 -688
rect -208 -689 -204 -668
rect -108 -689 -104 -668
rect -11 -689 -7 -635
rect 37 -649 41 -541
rect 212 -644 216 -435
rect 75 -648 216 -644
rect 37 -653 70 -649
rect 66 -680 70 -653
rect 75 -689 79 -648
rect -783 -793 -779 -692
rect -208 -693 -178 -689
rect -108 -693 -83 -689
rect -11 -693 6 -689
rect 75 -693 97 -689
rect -179 -714 164 -710
rect -744 -746 -635 -742
rect -744 -796 -740 -746
rect 148 -763 349 -759
rect -69 -776 -65 -769
rect -368 -780 -65 -776
rect -35 -778 94 -774
rect -368 -792 -364 -780
rect -35 -790 -31 -778
rect 90 -779 94 -778
rect 148 -779 152 -763
rect 90 -783 152 -779
rect 173 -790 179 -786
rect -124 -794 -31 -790
rect 175 -818 179 -790
rect 189 -811 193 -778
rect 189 -815 207 -811
rect 203 -818 207 -815
rect 232 -880 348 -876
rect 232 -881 236 -880
rect 218 -885 236 -881
rect 67 -956 97 -952
rect -1053 -962 -275 -958
rect -1053 -1189 -1049 -962
rect -1031 -970 -628 -966
rect -1031 -988 -1027 -970
rect -718 -993 -638 -989
rect -1053 -1193 -862 -1189
rect -866 -1584 -862 -1193
rect -789 -1317 -785 -1242
rect -718 -1287 -714 -993
rect -279 -994 -275 -962
rect 67 -963 71 -956
rect -229 -967 71 -963
rect -279 -998 -253 -994
rect 266 -1162 270 -1096
rect -695 -1188 -630 -1184
rect -654 -1261 -650 -1209
rect -634 -1253 -630 -1188
rect 392 -1191 396 -435
rect 185 -1195 396 -1191
rect -634 -1257 -432 -1253
rect -654 -1265 -453 -1261
rect -718 -1291 -482 -1287
rect -789 -1321 -512 -1317
rect -516 -1525 -512 -1321
rect -486 -1526 -482 -1291
rect -457 -1463 -453 -1265
rect -436 -1436 -432 -1257
rect -436 -1440 -351 -1436
rect -355 -1463 -351 -1440
rect -266 -1463 -262 -1315
rect 185 -1357 189 -1195
rect -182 -1361 189 -1357
rect -182 -1463 -178 -1361
rect -457 -1467 -414 -1463
rect -355 -1467 -332 -1463
rect -266 -1467 -243 -1463
rect -182 -1467 -159 -1463
rect -430 -1488 -415 -1484
rect -371 -1488 -333 -1484
rect -288 -1488 -244 -1484
rect -199 -1488 -160 -1484
rect -115 -1488 -98 -1484
rect -365 -1558 -361 -1519
rect -283 -1558 -279 -1519
rect -194 -1558 -190 -1519
rect -365 -1562 -160 -1558
rect -164 -1570 -160 -1562
rect -146 -1560 -142 -1547
rect -146 -1564 -2 -1560
rect -866 -1588 -16 -1584
rect -1001 -1602 -832 -1598
rect -1001 -1644 -997 -1602
rect -20 -1612 -16 -1588
rect -6 -1607 -2 -1564
rect -6 -1611 12 -1607
rect 8 -1614 12 -1611
rect -962 -1645 -958 -1631
rect -606 -1641 -602 -1622
rect -567 -1643 -563 -1621
rect -224 -1641 -220 -1631
rect -185 -1642 -181 -1631
rect -1244 -1846 -1230 -1842
rect -847 -1844 -836 -1840
rect -468 -1844 -455 -1840
rect -164 -1865 -160 -1829
rect -115 -1865 -111 -1858
rect -164 -1869 81 -1865
rect -1218 -2111 -1214 -2003
rect -820 -2111 -816 -2001
rect -1218 -2112 -816 -2111
rect -438 -2112 -434 -2001
rect -115 -2112 -111 -1869
rect -1218 -2115 -111 -2112
rect -818 -2116 -111 -2115
<< polycontact >>
rect 79 109 83 113
rect 0 88 4 92
rect 79 88 83 92
rect 162 88 166 92
rect 236 88 240 92
rect 71 55 75 59
rect 155 55 159 59
rect -606 -94 -601 -89
rect 57 23 61 28
rect 57 -23 61 -18
rect 138 23 142 28
rect 143 -23 147 -18
rect 221 23 225 28
rect 295 23 299 28
rect 227 -23 231 -18
rect 307 -23 311 -18
rect -445 -104 -441 -100
rect 57 -88 61 -83
rect -522 -125 -518 -121
rect -509 -137 -505 -132
rect -601 -242 -596 -237
rect -434 -114 -430 -109
rect -132 -113 -128 -109
rect -192 -155 -188 -151
rect -153 -157 -149 -153
rect -141 -163 -137 -158
rect -225 -333 -221 -329
rect -149 -333 -145 -329
rect -414 -370 -409 -366
rect -151 -416 -147 -412
rect 143 -88 147 -83
rect 227 -88 231 -83
rect 307 -88 311 -83
rect 125 -153 129 -149
rect -115 -158 -111 -154
rect 164 -155 168 -151
rect 299 -143 303 -139
rect 317 -142 321 -138
rect 225 -237 229 -232
rect -47 -356 -43 -352
rect -123 -503 -119 -499
rect 165 -414 170 -410
rect -123 -639 -119 -635
rect -695 -668 -691 -664
rect -440 -692 -436 -688
rect -7 -639 -3 -635
rect 66 -684 70 -680
rect -635 -746 -631 -742
rect 148 -759 152 -755
rect 349 -763 354 -759
rect -69 -769 -65 -764
rect -35 -774 -30 -769
rect 56 -774 61 -770
rect -407 -790 -403 -786
rect 189 -778 193 -773
rect 168 -790 173 -786
rect -129 -794 -124 -790
rect -22 -797 -18 -791
rect 17 -797 21 -793
rect 348 -880 352 -876
rect 214 -885 218 -881
rect 97 -956 101 -952
rect -628 -970 -624 -966
rect -1031 -992 -1027 -988
rect -1016 -999 -1012 -995
rect -742 -1057 -738 -1053
rect -789 -1242 -785 -1238
rect -233 -967 -229 -963
rect -366 -1051 -362 -1047
rect 19 -1056 23 -1052
rect 266 -1096 270 -1092
rect 266 -1166 270 -1162
rect -695 -1184 -691 -1180
rect -654 -1209 -650 -1205
rect -516 -1529 -512 -1525
rect -262 -1319 -258 -1315
rect -486 -1530 -482 -1526
rect -365 -1519 -361 -1515
rect -283 -1519 -279 -1515
rect -194 -1519 -190 -1515
rect -110 -1519 -106 -1515
rect -146 -1547 -142 -1543
rect -164 -1574 -160 -1570
rect -832 -1602 -828 -1598
rect -606 -1622 -602 -1618
rect -962 -1631 -958 -1627
rect -567 -1621 -563 -1617
rect -224 -1631 -220 -1627
rect -185 -1631 -181 -1627
rect -164 -1829 -160 -1825
rect -115 -1858 -111 -1854
rect 81 -1869 85 -1865
rect -960 -1904 -956 -1900
rect -565 -1902 -561 -1898
rect -183 -1902 -179 -1898
rect -1218 -2003 -1214 -1999
rect -820 -2001 -816 -1997
rect -438 -2001 -434 -1997
<< metal1 >>
rect -581 169 439 224
rect 58 124 63 169
rect 66 168 71 169
rect -58 119 63 124
rect 67 126 71 168
rect 67 122 447 126
rect -58 -77 -53 119
rect 67 115 71 122
rect -666 -82 -53 -77
rect -46 111 71 115
rect 79 113 437 117
rect -666 -655 -661 -82
rect -46 -85 -42 111
rect -140 -89 -42 -85
rect -37 98 75 102
rect -601 -93 -136 -89
rect -37 -93 -33 98
rect 71 59 75 98
rect 155 98 350 102
rect 155 59 159 98
rect 0 -26 6 28
rect 23 -7 27 5
rect 23 -12 77 -7
rect -601 -94 -430 -93
rect -794 -660 -661 -655
rect -654 -104 -445 -100
rect -794 -781 -789 -660
rect -1028 -786 -789 -781
rect -1028 -951 -1023 -786
rect -1063 -956 -1023 -951
rect -1063 -988 -1058 -956
rect -1063 -992 -1031 -988
rect -1027 -992 -994 -988
rect -1030 -999 -1016 -995
rect -1030 -1173 -1026 -999
rect -738 -1057 -702 -1053
rect -1030 -1177 -848 -1173
rect -852 -1618 -848 -1177
rect -748 -1274 -744 -1206
rect -708 -1246 -702 -1057
rect -695 -1180 -691 -668
rect -654 -1205 -650 -104
rect -434 -109 -430 -94
rect -132 -97 -33 -93
rect -132 -109 -128 -97
rect 21 -121 25 -106
rect -518 -125 25 -121
rect 72 -129 77 -12
rect 84 -25 90 29
rect 102 -9 106 5
rect 102 -13 155 -9
rect 88 -26 90 -25
rect -505 -137 -438 -132
rect -635 -182 -586 -178
rect -635 -742 -631 -182
rect -464 -298 -449 -294
rect -525 -350 -457 -343
rect -464 -713 -457 -350
rect -453 -620 -449 -298
rect -444 -515 -438 -137
rect -192 -133 77 -129
rect -192 -151 -188 -133
rect 106 -137 112 -106
rect 151 -126 155 -13
rect 168 -25 174 29
rect 185 -9 189 5
rect 236 -3 240 28
rect 236 -6 252 -3
rect 259 -4 263 4
rect 185 -13 243 -9
rect 172 -26 174 -25
rect -153 -142 112 -137
rect 125 -130 155 -126
rect 192 -130 196 -106
rect -153 -153 -149 -142
rect 125 -149 129 -130
rect 164 -134 196 -130
rect 238 -130 243 -13
rect 248 -24 252 -6
rect 271 -119 275 -106
rect 271 -123 321 -119
rect 164 -151 168 -134
rect 238 -135 303 -130
rect 299 -139 303 -135
rect 317 -138 321 -123
rect 346 -122 350 98
rect 346 -126 389 -122
rect -137 -163 -111 -158
rect -364 -333 -225 -329
rect -145 -333 -119 -329
rect -364 -360 -360 -333
rect -147 -416 -126 -412
rect -444 -520 -245 -515
rect -250 -607 -245 -520
rect -131 -521 -126 -416
rect -123 -499 -119 -333
rect -116 -345 -111 -163
rect 187 -182 234 -178
rect -116 -350 -92 -345
rect -47 -357 -43 -356
rect 187 -410 192 -182
rect 300 -349 340 -344
rect 170 -414 192 -410
rect 356 -413 360 -297
rect 195 -417 360 -413
rect 157 -421 199 -417
rect 385 -422 389 -126
rect 202 -426 389 -422
rect -131 -527 64 -521
rect -197 -607 -193 -591
rect -250 -612 -193 -607
rect -157 -620 -153 -564
rect 57 -607 64 -527
rect 119 -607 124 -589
rect 57 -612 124 -607
rect 160 -620 164 -563
rect -453 -624 164 -620
rect -187 -681 -183 -624
rect -123 -643 -111 -639
rect -436 -692 -378 -688
rect -464 -717 -403 -713
rect -407 -786 -403 -717
rect -382 -772 -378 -692
rect -163 -765 -159 -764
rect -164 -769 -159 -765
rect -163 -772 -159 -769
rect -382 -776 -159 -772
rect -129 -790 -124 -741
rect -115 -785 -111 -643
rect -92 -663 -88 -624
rect 202 -635 206 -426
rect -3 -639 322 -635
rect -92 -667 269 -663
rect -92 -683 -88 -667
rect -2 -682 2 -667
rect 89 -684 93 -667
rect -34 -741 -29 -736
rect -35 -769 -30 -741
rect 22 -782 26 -767
rect 56 -770 61 -741
rect -115 -789 -18 -785
rect -22 -791 -18 -789
rect 17 -786 26 -782
rect 66 -786 70 -684
rect 148 -755 152 -741
rect 112 -773 117 -764
rect 112 -778 189 -773
rect 17 -793 21 -786
rect 66 -790 168 -786
rect 48 -838 109 -834
rect -362 -1051 -341 -1047
rect -414 -1227 -408 -1226
rect -414 -1233 -407 -1227
rect -414 -1246 -408 -1233
rect -708 -1252 -408 -1246
rect -372 -1274 -368 -1200
rect -345 -1249 -341 -1051
rect 48 -1052 52 -838
rect 265 -950 269 -667
rect 232 -954 270 -950
rect 174 -1005 232 -1000
rect 175 -1006 180 -1005
rect 23 -1056 52 -1052
rect 266 -1088 270 -954
rect 68 -1092 270 -1088
rect -26 -1249 -22 -1233
rect -345 -1253 -22 -1249
rect 13 -1274 17 -1205
rect 68 -1274 72 -1092
rect 318 -1130 322 -639
rect 433 -710 437 113
rect -748 -1278 72 -1274
rect 113 -1134 322 -1130
rect 339 -714 437 -710
rect 113 -1315 117 -1134
rect -258 -1319 117 -1315
rect 266 -1172 270 -1166
rect 339 -1172 343 -714
rect 443 -759 447 122
rect 354 -763 447 -759
rect 414 -876 418 -763
rect 352 -880 418 -876
rect 266 -1176 343 -1172
rect 266 -1396 270 -1176
rect 414 -1224 418 -880
rect 49 -1400 270 -1396
rect 299 -1228 418 -1224
rect 49 -1427 53 -1400
rect 299 -1423 303 -1228
rect -424 -1431 53 -1427
rect -424 -1459 -420 -1431
rect -342 -1455 -338 -1431
rect -252 -1457 -248 -1431
rect -169 -1457 -165 -1431
rect -249 -1458 -248 -1457
rect -589 -1487 -441 -1483
rect -589 -1598 -585 -1487
rect -568 -1507 -460 -1503
rect -828 -1602 -585 -1598
rect -567 -1617 -563 -1507
rect -852 -1622 -606 -1618
rect -516 -1627 -512 -1529
rect -486 -1597 -482 -1530
rect -464 -1569 -460 -1507
rect -445 -1557 -441 -1487
rect -401 -1557 -397 -1539
rect -445 -1561 -397 -1557
rect -319 -1569 -315 -1538
rect -464 -1573 -315 -1569
rect -229 -1572 -225 -1538
rect -229 -1576 -181 -1572
rect -486 -1601 -220 -1597
rect -958 -1631 -512 -1627
rect -224 -1627 -220 -1601
rect -185 -1627 -181 -1576
rect -110 -1574 -106 -1519
rect -164 -1578 -106 -1574
rect -164 -1825 -160 -1578
rect -141 -1634 -86 -1630
rect -141 -1898 -137 -1634
rect 49 -1696 53 -1431
rect 81 -1427 303 -1423
rect 30 -1700 54 -1696
rect -21 -1801 26 -1796
rect -956 -1904 -926 -1900
rect -561 -1902 -532 -1898
rect -179 -1902 -137 -1898
rect -1218 -1999 -1213 -1994
rect -930 -2012 -926 -1904
rect -930 -2016 -672 -2012
rect -1007 -2093 -1002 -2083
rect -966 -2147 -962 -2053
rect -676 -2097 -672 -2016
rect -612 -2097 -608 -2082
rect -676 -2101 -608 -2097
rect -571 -2147 -567 -2050
rect -536 -2109 -532 -1902
rect -233 -2083 -223 -2077
rect -230 -2109 -226 -2083
rect -536 -2113 -226 -2109
rect -191 -2147 -187 -2050
rect -966 -2148 -187 -2147
rect 50 -2148 54 -1700
rect 81 -1865 85 -1427
rect -966 -2205 54 -2148
use full_adder  full_adder_7
timestamp 1669380902
transform 0 -1 -968 -1 0 -1646
box -7 -21 445 266
use full_adder  full_adder_6
timestamp 1669380902
transform 0 -1 -573 -1 0 -1644
box -7 -21 445 266
use full_adder  full_adder_5
timestamp 1669380902
transform 0 -1 -191 -1 0 -1644
box -7 -21 445 266
use half_adder  half_adder_3
timestamp 1669380902
transform -1 0 30 0 -1 -1812
box -11 -212 145 48
use full_adder  full_adder_4
timestamp 1669380902
transform 0 -1 -750 -1 0 -799
box -7 -21 445 266
use full_adder  full_adder_3
timestamp 1669380902
transform 0 -1 -374 -1 0 -793
box -7 -21 445 266
use edit  and_12
timestamp 1669377468
transform 0 1 -386 -1 0 -1455
box -6 -38 94 25
use edit  and_13
timestamp 1669377468
transform 0 1 -304 -1 0 -1455
box -6 -38 94 25
use edit  and_14
timestamp 1669377468
transform 0 1 -215 -1 0 -1455
box -6 -38 94 25
use edit  and_15
timestamp 1669377468
transform 0 1 -131 -1 0 -1455
box -6 -38 94 25
use full_adder  full_adder_2
timestamp 1669380902
transform 0 -1 11 -1 0 -798
box -7 -21 445 266
use edit  and_10
timestamp 1669377468
transform 0 1 36 -1 0 -681
box -6 -38 94 25
use edit  and_9
timestamp 1669377468
transform 0 1 -54 -1 0 -681
box -6 -38 94 25
use edit  and_8
timestamp 1669377468
transform 0 1 -149 -1 0 -681
box -6 -38 94 25
use edit  and_11
timestamp 1669377468
transform 0 1 127 -1 0 -681
box -6 -38 94 25
use half_adder  half_adder_2
timestamp 1669380902
transform -1 0 225 0 -1 -1016
box -11 -212 145 48
use half_adder  half_adder_1
timestamp 1669380902
transform -1 0 -472 0 -1 -360
box -11 -212 145 48
use full_adder  full_adder_1
timestamp 1669380902
transform 0 -1 -159 -1 0 -158
box -7 -21 445 266
use full_adder  full_adder_0
timestamp 1669380902
transform 0 -1 158 -1 0 -156
box -7 -21 445 266
use half_adder  half_adder_0
timestamp 1669380902
transform -1 0 349 0 -1 -360
box -11 -212 145 48
use edit  and_4
timestamp 1669377468
transform 0 1 36 -1 0 -23
box -6 -38 94 25
use edit  and_0
timestamp 1669377468
transform 0 1 38 -1 0 88
box -6 -38 94 25
use edit  and_7
timestamp 1669377468
transform 0 1 286 -1 0 -23
box -6 -38 94 25
use edit  and_6
timestamp 1669377468
transform 0 1 206 -1 0 -23
box -6 -38 94 25
use edit  and_3
timestamp 1669377468
transform 0 1 274 -1 0 88
box -6 -38 94 25
use edit  and_2
timestamp 1669377468
transform 0 1 200 -1 0 88
box -6 -38 94 25
use edit  and_5
timestamp 1669377468
transform 0 1 122 -1 0 -23
box -6 -38 94 25
use edit  and_1
timestamp 1669377468
transform 0 1 117 -1 0 88
box -6 -38 94 25
<< labels >>
rlabel polysilicon -5 57 -5 57 3 a3
rlabel polysilicon 309 78 309 78 7 b0
rlabel polysilicon 233 57 233 57 1 a0
rlabel polysilicon 316 -54 316 -54 7 b1
rlabel polysilicon 73 49 73 49 1 a2
rlabel polysilicon 157 53 157 53 1 a1
rlabel polysilicon 161 -712 161 -712 1 b2
rlabel polysilicon -102 -1486 -102 -1486 1 b3
rlabel metal1 -145 195 -145 195 1 vdd
rlabel metal1 -541 -2176 -541 -2176 1 gnd
rlabel metal1 261 -2 261 -2 1 p0
rlabel metal1 335 -347 335 -347 1 p1
rlabel metal1 224 -1002 224 -1002 1 p2
rlabel metal1 21 -1799 21 -1799 1 p3
rlabel polysilicon -463 -1842 -463 -1842 1 p4
rlabel polysilicon -841 -1842 -841 -1842 1 p5
rlabel polysilicon -1237 -1844 -1237 -1844 1 p6
rlabel metal1 -1005 -2090 -1005 -2090 1 p7
<< end >>
