AND2 MAGIC CIRCUIT 


.include TSMC_180nm.txt
.global gnd vdd
.option scale=0.01u

*********
*netlist*
*********

Vdd vdd gnd 1

M1000 out a_19_7# gnd Gnd CMOSN w=36 l=36
+  ad=5184 pd=360 as=12636 ps=738
M1001 vdd b a_19_7# vdd CMOSP w=144 l=36
+  ad=38232 pd=1422 as=24624 ps=630
M1002 a_19_7# b a_19_n19# Gnd CMOSN w=72 l=36
+  ad=6480 pd=324 as=12312 ps=486
M1003 a_19_n19# a gnd Gnd CMOSN w=72 l=36
+  ad=0 pd=0 as=0 ps=0
M1004 out a_19_7# vdd vdd CMOSP w=72 l=36
+  ad=10368 pd=432 as=0 ps=0
M1005 a_19_7# a vdd vdd CMOSP w=144 l=36
+  ad=0 pd=0 as=0 ps=0
C0 w_64_0# Gnd 1.51fF
C1 w_n1_0# Gnd 1.72fF

cout out gnd 10f

Va a gnd pulse(0 1 0 0.1u 0.1u 10u 20u)
Vb b gnd pulse(0 1 0 0.1u 0.1u 20u 40u) 


*control*
.control
tran 0.1u 100u

plot v(out) 
plot   v(a)
plot   v(b)

let delay_and_lh = 0
let delay_and_hl = 0

meas tran delay_and_lh trig v(a) val = 0.5 rise = 1 targ v(out) val = 0.5 rise = 1
meas tran delay_and_hl trig v(a) val = 0.5 fall = 1 targ v(out) val = 0.5 fall = 1
let prop_del_and = (delay_and_lh + -1*delay_and_hl)/2

echo                                              " ---------------------------------"  > "and_delays.txt"
echo 				   	  "|-> low to high delay = " "$&delay_and_lh|" >> "and_delays.txt"
echo 					  "|-> high to low delay = " "$&delay_and_hl|" >> "and_delays.txt"
echo "|-> average propogation delay = "                              "$&prop_del_and|" >> "and_delays.txt"
echo                             		  " ---------------------------------" >> "and_delays.txt"

.endc

.end
